
module Shifter( dataA, dataB, dataOut );
  input [31:0] dataA ;
  input [4:0] dataB ;
  output [31:0] dataOut ;

  wire [31:0] temp_1, temp_2, temp_4, temp_8, temp_16, temp ;


  assign temp_1[0] = ( dataB[0] ) ? 1'b0     : dataA[0] ;
  assign temp_1[1] = ( dataB[0] ) ? dataA[0] : dataA[1] ;
  assign temp_1[2] = ( dataB[0] ) ? dataA[1] : dataA[2] ;
  assign temp_1[3] = ( dataB[0] ) ? dataA[2] : dataA[3] ;
  assign temp_1[4] = ( dataB[0] ) ? dataA[3] : dataA[4] ;
  assign temp_1[5] = ( dataB[0] ) ? dataA[4] : dataA[5] ;
  assign temp_1[6] = ( dataB[0] ) ? dataA[5] : dataA[6] ;
  assign temp_1[7] = ( dataB[0] ) ? dataA[6] : dataA[7] ;
  assign temp_1[8] = ( dataB[0] ) ? dataA[7] : dataA[8] ;
  assign temp_1[9] = ( dataB[0] ) ? dataA[8] : dataA[9] ;
  assign temp_1[10] = ( dataB[0] ) ? dataA[9] : dataA[10] ;
  assign temp_1[11] = ( dataB[0] ) ? dataA[10] : dataA[11] ;
  assign temp_1[12] = ( dataB[0] ) ? dataA[11] : dataA[12] ;
  assign temp_1[13] = ( dataB[0] ) ? dataA[12] : dataA[13] ;
  assign temp_1[14] = ( dataB[0] ) ? dataA[13] : dataA[14] ;
  assign temp_1[15] = ( dataB[0] ) ? dataA[14] : dataA[15] ;
  assign temp_1[16] = ( dataB[0] ) ? dataA[15] : dataA[16] ;
  assign temp_1[17] = ( dataB[0] ) ? dataA[16] : dataA[17] ;
  assign temp_1[18] = ( dataB[0] ) ? dataA[17] : dataA[18] ;
  assign temp_1[19] = ( dataB[0] ) ? dataA[18] : dataA[19] ;
  assign temp_1[20] = ( dataB[0] ) ? dataA[19] : dataA[20] ;
  assign temp_1[21] = ( dataB[0] ) ? dataA[20] : dataA[21] ;
  assign temp_1[22] = ( dataB[0] ) ? dataA[21] : dataA[22] ;
  assign temp_1[23] = ( dataB[0] ) ? dataA[22] : dataA[23] ;
  assign temp_1[24] = ( dataB[0] ) ? dataA[23] : dataA[24] ;
  assign temp_1[25] = ( dataB[0] ) ? dataA[24] : dataA[25] ;
  assign temp_1[26] = ( dataB[0] ) ? dataA[25] : dataA[26] ;
  assign temp_1[27] = ( dataB[0] ) ? dataA[26] : dataA[27] ;
  assign temp_1[28] = ( dataB[0] ) ? dataA[27] : dataA[28] ;
  assign temp_1[29] = ( dataB[0] ) ? dataA[28] : dataA[29] ;
  assign temp_1[30] = ( dataB[0] ) ? dataA[29] : dataA[30] ;
  assign temp_1[31] = ( dataB[0] ) ? dataA[30] : dataA[31] ;


  assign temp_2[0] = ( dataB[1] ) ? 1'b0      : temp_1[0];
  assign temp_2[1] = ( dataB[1] ) ? 1'b0      : temp_1[1];
  assign temp_2[2] = ( dataB[1] ) ? temp_1[0] : temp_1[2] ;
  assign temp_2[3] = ( dataB[1] ) ? temp_1[1] : temp_1[3] ;
  assign temp_2[4] = ( dataB[1] ) ? temp_1[2] : temp_1[4] ;
  assign temp_2[5] = ( dataB[1] ) ? temp_1[3] : temp_1[5] ;
  assign temp_2[6] = ( dataB[1] ) ? temp_1[4] : temp_1[6] ;
  assign temp_2[7] = ( dataB[1] ) ? temp_1[5] : temp_1[7] ;
  assign temp_2[8] = ( dataB[1] ) ? temp_1[6] : temp_1[8] ;
  assign temp_2[9] = ( dataB[1] ) ? temp_1[7] : temp_1[9] ;
  assign temp_2[10] = ( dataB[1] ) ? temp_1[8] : temp_1[10] ;
  assign temp_2[11] = ( dataB[1] ) ? temp_1[9] : temp_1[11] ;
  assign temp_2[12] = ( dataB[1] ) ? temp_1[10] : temp_1[12] ;
  assign temp_2[13] = ( dataB[1] ) ? temp_1[11] : temp_1[13] ;
  assign temp_2[14] = ( dataB[1] ) ? temp_1[12] : temp_1[14] ;
  assign temp_2[15] = ( dataB[1] ) ? temp_1[13] : temp_1[15] ;
  assign temp_2[16] = ( dataB[1] ) ? temp_1[14] : temp_1[16] ;
  assign temp_2[17] = ( dataB[1] ) ? temp_1[15] : temp_1[17] ;
  assign temp_2[18] = ( dataB[1] ) ? temp_1[16] : temp_1[18] ;
  assign temp_2[19] = ( dataB[1] ) ? temp_1[17] : temp_1[19] ;
  assign temp_2[20] = ( dataB[1] ) ? temp_1[18] : temp_1[20] ;
  assign temp_2[21] = ( dataB[1] ) ? temp_1[19] : temp_1[21] ;
  assign temp_2[22] = ( dataB[1] ) ? temp_1[20] : temp_1[22] ;
  assign temp_2[23] = ( dataB[1] ) ? temp_1[21] : temp_1[23] ;
  assign temp_2[24] = ( dataB[1] ) ? temp_1[22] : temp_1[24] ;
  assign temp_2[25] = ( dataB[1] ) ? temp_1[23] : temp_1[25] ;
  assign temp_2[26] = ( dataB[1] ) ? temp_1[24] : temp_1[26] ;
  assign temp_2[27] = ( dataB[1] ) ? temp_1[25] : temp_1[27] ;
  assign temp_2[28] = ( dataB[1] ) ? temp_1[26] : temp_1[28] ;
  assign temp_2[29] = ( dataB[1] ) ? temp_1[27] : temp_1[29] ;
  assign temp_2[30] = ( dataB[1] ) ? temp_1[28] : temp_1[30] ;
  assign temp_2[31] = ( dataB[1] ) ? temp_1[29] : temp_1[31] ;


  assign temp_4[0] = ( dataB[2] ) ? 1'b0      : temp_2[0] ;
  assign temp_4[1] = ( dataB[2] ) ? 1'b0      : temp_2[1] ;
  assign temp_4[2] = ( dataB[2] ) ? 1'b0      : temp_2[2] ;
  assign temp_4[3] = ( dataB[2] ) ? 1'b0      : temp_2[3] ;
  assign temp_4[4] = ( dataB[2] ) ? temp_2[0] : temp_2[4] ;
  assign temp_4[5] = ( dataB[2] ) ? temp_2[1] : temp_2[5] ;
  assign temp_4[6] = ( dataB[2] ) ? temp_2[2] : temp_2[6] ;
  assign temp_4[7] = ( dataB[2] ) ? temp_2[3] : temp_2[7] ;
  assign temp_4[8] = ( dataB[2] ) ? temp_2[4] : temp_2[8] ;
  assign temp_4[9] = ( dataB[2] ) ? temp_2[5] : temp_2[9] ;
  assign temp_4[10] = ( dataB[2] ) ? temp_2[6] : temp_2[10] ;
  assign temp_4[11] = ( dataB[2] ) ? temp_2[7] : temp_2[11] ;
  assign temp_4[12] = ( dataB[2] ) ? temp_2[8] : temp_2[12] ;
  assign temp_4[13] = ( dataB[2] ) ? temp_2[9] : temp_2[13] ;
  assign temp_4[14] = ( dataB[2] ) ? temp_2[10] : temp_2[14] ;
  assign temp_4[15] = ( dataB[2] ) ? temp_2[11] : temp_2[15] ;
  assign temp_4[16] = ( dataB[2] ) ? temp_2[12] : temp_2[16] ;
  assign temp_4[17] = ( dataB[2] ) ? temp_2[13] : temp_2[17] ;
  assign temp_4[18] = ( dataB[2] ) ? temp_2[14] : temp_2[18] ;
  assign temp_4[19] = ( dataB[2] ) ? temp_2[15] : temp_2[19] ;
  assign temp_4[20] = ( dataB[2] ) ? temp_2[16] : temp_2[20] ;
  assign temp_4[21] = ( dataB[2] ) ? temp_2[17] : temp_2[21] ;
  assign temp_4[22] = ( dataB[2] ) ? temp_2[18] : temp_2[22] ;
  assign temp_4[23] = ( dataB[2] ) ? temp_2[19] : temp_2[23] ;
  assign temp_4[24] = ( dataB[2] ) ? temp_2[20] : temp_2[24] ;
  assign temp_4[25] = ( dataB[2] ) ? temp_2[21] : temp_2[25] ;
  assign temp_4[26] = ( dataB[2] ) ? temp_2[22] : temp_2[26] ;
  assign temp_4[27] = ( dataB[2] ) ? temp_2[23] : temp_2[27] ;
  assign temp_4[28] = ( dataB[2] ) ? temp_2[24] : temp_2[28] ;
  assign temp_4[29] = ( dataB[2] ) ? temp_2[25] : temp_2[29] ;
  assign temp_4[30] = ( dataB[2] ) ? temp_2[26] : temp_2[30] ;
  assign temp_4[31] = ( dataB[2] ) ? temp_2[27] : temp_2[31] ;


  assign temp_8[0] = ( dataB[3] ) ? 1'b0      : temp_4[0] ;
  assign temp_8[1] = ( dataB[3] ) ? 1'b0      : temp_4[1] ;
  assign temp_8[2] = ( dataB[3] ) ? 1'b0      : temp_4[2] ;
  assign temp_8[3] = ( dataB[3] ) ? 1'b0      : temp_4[3] ;
  assign temp_8[4] = ( dataB[3] ) ? 1'b0      : temp_4[4] ;
  assign temp_8[5] = ( dataB[3] ) ? 1'b0      : temp_4[5] ;
  assign temp_8[6] = ( dataB[3] ) ? 1'b0      : temp_4[6] ;
  assign temp_8[7] = ( dataB[3] ) ? 1'b0      : temp_4[7] ;
  assign temp_8[8] = ( dataB[3] ) ? temp_4[0] : temp_4[8] ;
  assign temp_8[9] = ( dataB[3] ) ? temp_4[1] : temp_4[9] ;
  assign temp_8[10] = ( dataB[3] ) ? temp_4[2] : temp_4[10] ;
  assign temp_8[11] = ( dataB[3] ) ? temp_4[3] : temp_4[11] ;
  assign temp_8[12] = ( dataB[3] ) ? temp_4[4] : temp_4[12] ;
  assign temp_8[13] = ( dataB[3] ) ? temp_4[5] : temp_4[13] ;
  assign temp_8[14] = ( dataB[3] ) ? temp_4[6] : temp_4[14] ;
  assign temp_8[15] = ( dataB[3] ) ? temp_4[7] : temp_4[15] ;
  assign temp_8[16] = ( dataB[3] ) ? temp_4[8] : temp_4[16] ;
  assign temp_8[17] = ( dataB[3] ) ? temp_4[9] : temp_4[17] ;
  assign temp_8[18] = ( dataB[3] ) ? temp_4[10] : temp_4[18] ;
  assign temp_8[19] = ( dataB[3] ) ? temp_4[11] : temp_4[19] ;
  assign temp_8[20] = ( dataB[3] ) ? temp_4[12] : temp_4[20] ;
  assign temp_8[21] = ( dataB[3] ) ? temp_4[13] : temp_4[21] ;
  assign temp_8[22] = ( dataB[3] ) ? temp_4[14] : temp_4[22] ;
  assign temp_8[23] = ( dataB[3] ) ? temp_4[15] : temp_4[23] ;
  assign temp_8[24] = ( dataB[3] ) ? temp_4[16] : temp_4[24] ;
  assign temp_8[25] = ( dataB[3] ) ? temp_4[17] : temp_4[25] ;
  assign temp_8[26] = ( dataB[3] ) ? temp_4[18] : temp_4[26] ;
  assign temp_8[27] = ( dataB[3] ) ? temp_4[19] : temp_4[27] ;
  assign temp_8[28] = ( dataB[3] ) ? temp_4[20] : temp_4[28] ;
  assign temp_8[29] = ( dataB[3] ) ? temp_4[21] : temp_4[29] ;
  assign temp_8[30] = ( dataB[3] ) ? temp_4[22] : temp_4[30] ;
  assign temp_8[31] = ( dataB[3] ) ? temp_4[23] : temp_4[31] ;


  assign temp_16[0] = ( dataB[4] ) ? 1'b0      : temp_8[0] ;
  assign temp_16[1] = ( dataB[4] ) ? 1'b0      : temp_8[1] ;
  assign temp_16[2] = ( dataB[4] ) ? 1'b0      : temp_8[2] ;
  assign temp_16[3] = ( dataB[4] ) ? 1'b0      : temp_8[3] ;
  assign temp_16[4] = ( dataB[4] ) ? 1'b0      : temp_8[4] ;
  assign temp_16[5] = ( dataB[4] ) ? 1'b0      : temp_8[5] ;
  assign temp_16[6] = ( dataB[4] ) ? 1'b0      : temp_8[6] ;
  assign temp_16[7] = ( dataB[4] ) ? 1'b0      : temp_8[7] ;
  assign temp_16[8] = ( dataB[4] ) ? 1'b0      : temp_8[8] ;
  assign temp_16[9] = ( dataB[4] ) ? 1'b0      : temp_8[9] ;
  assign temp_16[10] = ( dataB[4] ) ? 1'b0      : temp_8[10] ;
  assign temp_16[11] = ( dataB[4] ) ? 1'b0      : temp_8[11] ;
  assign temp_16[12] = ( dataB[4] ) ? 1'b0      : temp_8[12] ;
  assign temp_16[13] = ( dataB[4] ) ? 1'b0      : temp_8[13] ;
  assign temp_16[14] = ( dataB[4] ) ? 1'b0      : temp_8[14] ;
  assign temp_16[15] = ( dataB[4] ) ? 1'b0      : temp_8[15] ;
  assign temp_16[16] = ( dataB[4] ) ? temp_8[0] : temp_8[16] ;
  assign temp_16[17] = ( dataB[4] ) ? temp_8[1] : temp_8[17] ;
  assign temp_16[18] = ( dataB[4] ) ? temp_8[2] : temp_8[18] ;
  assign temp_16[19] = ( dataB[4] ) ? temp_8[3] : temp_8[19] ;
  assign temp_16[20] = ( dataB[4] ) ? temp_8[4] : temp_8[20] ;
  assign temp_16[21] = ( dataB[4] ) ? temp_8[5] : temp_8[21] ;
  assign temp_16[22] = ( dataB[4] ) ? temp_8[6] : temp_8[22] ;
  assign temp_16[23] = ( dataB[4] ) ? temp_8[7] : temp_8[23] ;
  assign temp_16[24] = ( dataB[4] ) ? temp_8[8] : temp_8[24] ;
  assign temp_16[25] = ( dataB[4] ) ? temp_8[9] : temp_8[25] ;
  assign temp_16[26] = ( dataB[4] ) ? temp_8[10] : temp_8[26] ;
  assign temp_16[27] = ( dataB[4] ) ? temp_8[11] : temp_8[27] ;
  assign temp_16[28] = ( dataB[4] ) ? temp_8[12] : temp_8[28] ;
  assign temp_16[29] = ( dataB[4] ) ? temp_8[13] : temp_8[29] ;
  assign temp_16[30] = ( dataB[4] ) ? temp_8[14] : temp_8[30] ;
  assign temp_16[31] = ( dataB[4] ) ? temp_8[15] : temp_8[31] ;

  assign temp = temp_16 ;
  assign dataOut = temp ;

endmodule
